library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

PACKAGE BUFFON2 IS
type padded_arrray_t is array (0 to 63) of std_logic_vector(511 downto 0) ;
END PACKAGE BUFFON2;